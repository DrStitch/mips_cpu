`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/02/22 16:02:31
// Design Name: 
// Module Name: MEM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MEM(
	in_pc,
	in_ir,
	in_signal,
	in_dst,
	in_r2,
	in_r,
	in_v0,
	in_a0
    out_pc,
    out_ir,
    out_signal,
    out_dst,
    out_d,
    out_r,
    out_v0,
    out_a0
    );
endmodule
